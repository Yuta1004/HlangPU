action_table[0] = 10'h1_09; action_table[1] = 10'h1_03; action_table[2] = 10'h1_04; action_table[3] = 10'h0_00; action_table[4] = 10'h1_05; action_table[5] = 10'h1_06; action_table[6] = 10'h1_07; action_table[7] = 10'h1_0a; action_table[8] = 10'h0_00; action_table[9] = 10'h0_00; action_table[10] = 10'h0_00; action_table[11] = 10'h0_00; action_table[12] = 10'h0_00; action_table[13] = 10'h0_00; action_table[14] = 10'h0_00; action_table[15] = 10'h0_00;
action_table[16] = 10'h1_09; action_table[17] = 10'h1_03; action_table[18] = 10'h1_04; action_table[19] = 10'h0_00; action_table[20] = 10'h1_05; action_table[21] = 10'h1_06; action_table[22] = 10'h1_07; action_table[23] = 10'h1_0a; action_table[24] = 10'h0_00; action_table[25] = 10'h0_00; action_table[26] = 10'h0_00; action_table[27] = 10'h0_00; action_table[28] = 10'h2_01; action_table[29] = 10'h0_00; action_table[30] = 10'h0_00; action_table[31] = 10'h0_00;
action_table[32] = 10'h0_00; action_table[33] = 10'h0_00; action_table[34] = 10'h0_00; action_table[35] = 10'h0_00; action_table[36] = 10'h0_00; action_table[37] = 10'h0_00; action_table[38] = 10'h0_00; action_table[39] = 10'h0_00; action_table[40] = 10'h0_00; action_table[41] = 10'h1_0d; action_table[42] = 10'h1_0e; action_table[43] = 10'h1_0c; action_table[44] = 10'h0_00; action_table[45] = 10'h0_00; action_table[46] = 10'h0_00; action_table[47] = 10'h0_00;
action_table[48] = 10'h1_09; action_table[49] = 10'h0_00; action_table[50] = 10'h0_00; action_table[51] = 10'h0_00; action_table[52] = 10'h0_00; action_table[53] = 10'h0_00; action_table[54] = 10'h0_00; action_table[55] = 10'h1_0a; action_table[56] = 10'h0_00; action_table[57] = 10'h0_00; action_table[58] = 10'h0_00; action_table[59] = 10'h0_00; action_table[60] = 10'h0_00; action_table[61] = 10'h0_00; action_table[62] = 10'h0_00; action_table[63] = 10'h0_00;
action_table[64] = 10'h0_00; action_table[65] = 10'h0_00; action_table[66] = 10'h0_00; action_table[67] = 10'h1_10; action_table[68] = 10'h0_00; action_table[69] = 10'h0_00; action_table[70] = 10'h0_00; action_table[71] = 10'h0_00; action_table[72] = 10'h0_00; action_table[73] = 10'h0_00; action_table[74] = 10'h0_00; action_table[75] = 10'h0_00; action_table[76] = 10'h0_00; action_table[77] = 10'h0_00; action_table[78] = 10'h0_00; action_table[79] = 10'h0_00;
action_table[80] = 10'h0_00; action_table[81] = 10'h0_00; action_table[82] = 10'h0_00; action_table[83] = 10'h1_11; action_table[84] = 10'h0_00; action_table[85] = 10'h0_00; action_table[86] = 10'h0_00; action_table[87] = 10'h0_00; action_table[88] = 10'h0_00; action_table[89] = 10'h0_00; action_table[90] = 10'h0_00; action_table[91] = 10'h0_00; action_table[92] = 10'h0_00; action_table[93] = 10'h0_00; action_table[94] = 10'h0_00; action_table[95] = 10'h0_00;
action_table[96] = 10'h0_00; action_table[97] = 10'h0_00; action_table[98] = 10'h0_00; action_table[99] = 10'h1_12; action_table[100] = 10'h0_00; action_table[101] = 10'h0_00; action_table[102] = 10'h0_00; action_table[103] = 10'h0_00; action_table[104] = 10'h0_00; action_table[105] = 10'h0_00; action_table[106] = 10'h0_00; action_table[107] = 10'h0_00; action_table[108] = 10'h0_00; action_table[109] = 10'h0_00; action_table[110] = 10'h0_00; action_table[111] = 10'h0_00;
action_table[112] = 10'h0_00; action_table[113] = 10'h0_00; action_table[114] = 10'h0_00; action_table[115] = 10'h0_00; action_table[116] = 10'h0_00; action_table[117] = 10'h0_00; action_table[118] = 10'h0_00; action_table[119] = 10'h1_13; action_table[120] = 10'h0_00; action_table[121] = 10'h0_00; action_table[122] = 10'h0_00; action_table[123] = 10'h0_00; action_table[124] = 10'h0_00; action_table[125] = 10'h0_00; action_table[126] = 10'h0_00; action_table[127] = 10'h0_00;
action_table[128] = 10'h0_00; action_table[129] = 10'h0_00; action_table[130] = 10'h0_00; action_table[131] = 10'h0_00; action_table[132] = 10'h0_00; action_table[133] = 10'h0_00; action_table[134] = 10'h0_00; action_table[135] = 10'h0_00; action_table[136] = 10'h0_00; action_table[137] = 10'h2_0a; action_table[138] = 10'h2_0a; action_table[139] = 10'h2_0a; action_table[140] = 10'h0_00; action_table[141] = 10'h0_00; action_table[142] = 10'h0_00; action_table[143] = 10'h0_00;
action_table[144] = 10'h0_00; action_table[145] = 10'h0_00; action_table[146] = 10'h0_00; action_table[147] = 10'h0_00; action_table[148] = 10'h0_00; action_table[149] = 10'h0_00; action_table[150] = 10'h0_00; action_table[151] = 10'h0_00; action_table[152] = 10'h0_00; action_table[153] = 10'h2_0b; action_table[154] = 10'h2_0b; action_table[155] = 10'h2_0b; action_table[156] = 10'h0_00; action_table[157] = 10'h0_00; action_table[158] = 10'h0_00; action_table[159] = 10'h0_00;
action_table[160] = 10'h1_16; action_table[161] = 10'h0_00; action_table[162] = 10'h0_00; action_table[163] = 10'h0_00; action_table[164] = 10'h0_00; action_table[165] = 10'h0_00; action_table[166] = 10'h0_00; action_table[167] = 10'h1_17; action_table[168] = 10'h0_00; action_table[169] = 10'h0_00; action_table[170] = 10'h0_00; action_table[171] = 10'h0_00; action_table[172] = 10'h0_00; action_table[173] = 10'h0_00; action_table[174] = 10'h0_00; action_table[175] = 10'h0_00;
action_table[176] = 10'h0_00; action_table[177] = 10'h0_00; action_table[178] = 10'h0_00; action_table[179] = 10'h0_00; action_table[180] = 10'h0_00; action_table[181] = 10'h0_00; action_table[182] = 10'h0_00; action_table[183] = 10'h0_00; action_table[184] = 10'h0_00; action_table[185] = 10'h0_00; action_table[186] = 10'h0_00; action_table[187] = 10'h0_00; action_table[188] = 10'h3_00; action_table[189] = 10'h0_00; action_table[190] = 10'h0_00; action_table[191] = 10'h0_00;
action_table[192] = 10'h2_02; action_table[193] = 10'h2_02; action_table[194] = 10'h2_02; action_table[195] = 10'h0_00; action_table[196] = 10'h2_02; action_table[197] = 10'h2_02; action_table[198] = 10'h2_02; action_table[199] = 10'h2_02; action_table[200] = 10'h0_00; action_table[201] = 10'h0_00; action_table[202] = 10'h0_00; action_table[203] = 10'h0_00; action_table[204] = 10'h2_02; action_table[205] = 10'h0_00; action_table[206] = 10'h0_00; action_table[207] = 10'h0_00;
action_table[208] = 10'h1_09; action_table[209] = 10'h0_00; action_table[210] = 10'h0_00; action_table[211] = 10'h0_00; action_table[212] = 10'h0_00; action_table[213] = 10'h0_00; action_table[214] = 10'h0_00; action_table[215] = 10'h1_0a; action_table[216] = 10'h0_00; action_table[217] = 10'h0_00; action_table[218] = 10'h0_00; action_table[219] = 10'h0_00; action_table[220] = 10'h0_00; action_table[221] = 10'h0_00; action_table[222] = 10'h0_00; action_table[223] = 10'h0_00;
action_table[224] = 10'h1_09; action_table[225] = 10'h0_00; action_table[226] = 10'h0_00; action_table[227] = 10'h0_00; action_table[228] = 10'h0_00; action_table[229] = 10'h0_00; action_table[230] = 10'h0_00; action_table[231] = 10'h1_0a; action_table[232] = 10'h0_00; action_table[233] = 10'h0_00; action_table[234] = 10'h0_00; action_table[235] = 10'h0_00; action_table[236] = 10'h0_00; action_table[237] = 10'h0_00; action_table[238] = 10'h0_00; action_table[239] = 10'h0_00;
action_table[240] = 10'h0_00; action_table[241] = 10'h0_00; action_table[242] = 10'h0_00; action_table[243] = 10'h0_00; action_table[244] = 10'h0_00; action_table[245] = 10'h0_00; action_table[246] = 10'h0_00; action_table[247] = 10'h0_00; action_table[248] = 10'h0_00; action_table[249] = 10'h1_0d; action_table[250] = 10'h1_0e; action_table[251] = 10'h1_1a; action_table[252] = 10'h0_00; action_table[253] = 10'h0_00; action_table[254] = 10'h0_00; action_table[255] = 10'h0_00;
action_table[256] = 10'h1_09; action_table[257] = 10'h0_00; action_table[258] = 10'h0_00; action_table[259] = 10'h0_00; action_table[260] = 10'h0_00; action_table[261] = 10'h0_00; action_table[262] = 10'h0_00; action_table[263] = 10'h1_0a; action_table[264] = 10'h0_00; action_table[265] = 10'h0_00; action_table[266] = 10'h0_00; action_table[267] = 10'h0_00; action_table[268] = 10'h0_00; action_table[269] = 10'h0_00; action_table[270] = 10'h0_00; action_table[271] = 10'h0_00;
action_table[272] = 10'h1_09; action_table[273] = 10'h0_00; action_table[274] = 10'h0_00; action_table[275] = 10'h0_00; action_table[276] = 10'h0_00; action_table[277] = 10'h0_00; action_table[278] = 10'h0_00; action_table[279] = 10'h1_0a; action_table[280] = 10'h0_00; action_table[281] = 10'h0_00; action_table[282] = 10'h0_00; action_table[283] = 10'h0_00; action_table[284] = 10'h0_00; action_table[285] = 10'h0_00; action_table[286] = 10'h0_00; action_table[287] = 10'h0_00;
action_table[288] = 10'h1_09; action_table[289] = 10'h0_00; action_table[290] = 10'h0_00; action_table[291] = 10'h0_00; action_table[292] = 10'h0_00; action_table[293] = 10'h0_00; action_table[294] = 10'h0_00; action_table[295] = 10'h1_0a; action_table[296] = 10'h0_00; action_table[297] = 10'h0_00; action_table[298] = 10'h0_00; action_table[299] = 10'h0_00; action_table[300] = 10'h0_00; action_table[301] = 10'h0_00; action_table[302] = 10'h0_00; action_table[303] = 10'h0_00;
action_table[304] = 10'h1_16; action_table[305] = 10'h0_00; action_table[306] = 10'h0_00; action_table[307] = 10'h0_00; action_table[308] = 10'h0_00; action_table[309] = 10'h0_00; action_table[310] = 10'h0_00; action_table[311] = 10'h1_17; action_table[312] = 10'h0_00; action_table[313] = 10'h0_00; action_table[314] = 10'h0_00; action_table[315] = 10'h0_00; action_table[316] = 10'h0_00; action_table[317] = 10'h0_00; action_table[318] = 10'h0_00; action_table[319] = 10'h0_00;
action_table[320] = 10'h0_00; action_table[321] = 10'h0_00; action_table[322] = 10'h0_00; action_table[323] = 10'h0_00; action_table[324] = 10'h0_00; action_table[325] = 10'h0_00; action_table[326] = 10'h0_00; action_table[327] = 10'h0_00; action_table[328] = 10'h1_1f; action_table[329] = 10'h1_20; action_table[330] = 10'h1_21; action_table[331] = 10'h0_00; action_table[332] = 10'h0_00; action_table[333] = 10'h0_00; action_table[334] = 10'h0_00; action_table[335] = 10'h0_00;
action_table[336] = 10'h0_00; action_table[337] = 10'h0_00; action_table[338] = 10'h0_00; action_table[339] = 10'h0_00; action_table[340] = 10'h0_00; action_table[341] = 10'h0_00; action_table[342] = 10'h0_00; action_table[343] = 10'h0_00; action_table[344] = 10'h2_0a; action_table[345] = 10'h2_0a; action_table[346] = 10'h2_0a; action_table[347] = 10'h0_00; action_table[348] = 10'h0_00; action_table[349] = 10'h0_00; action_table[350] = 10'h0_00; action_table[351] = 10'h0_00;
action_table[352] = 10'h0_00; action_table[353] = 10'h0_00; action_table[354] = 10'h0_00; action_table[355] = 10'h0_00; action_table[356] = 10'h0_00; action_table[357] = 10'h0_00; action_table[358] = 10'h0_00; action_table[359] = 10'h0_00; action_table[360] = 10'h2_0b; action_table[361] = 10'h2_0b; action_table[362] = 10'h2_0b; action_table[363] = 10'h0_00; action_table[364] = 10'h0_00; action_table[365] = 10'h0_00; action_table[366] = 10'h0_00; action_table[367] = 10'h0_00;
action_table[368] = 10'h1_16; action_table[369] = 10'h0_00; action_table[370] = 10'h0_00; action_table[371] = 10'h0_00; action_table[372] = 10'h0_00; action_table[373] = 10'h0_00; action_table[374] = 10'h0_00; action_table[375] = 10'h1_17; action_table[376] = 10'h0_00; action_table[377] = 10'h0_00; action_table[378] = 10'h0_00; action_table[379] = 10'h0_00; action_table[380] = 10'h0_00; action_table[381] = 10'h0_00; action_table[382] = 10'h0_00; action_table[383] = 10'h0_00;
action_table[384] = 10'h0_00; action_table[385] = 10'h0_00; action_table[386] = 10'h0_00; action_table[387] = 10'h0_00; action_table[388] = 10'h0_00; action_table[389] = 10'h0_00; action_table[390] = 10'h0_00; action_table[391] = 10'h0_00; action_table[392] = 10'h0_00; action_table[393] = 10'h2_08; action_table[394] = 10'h2_08; action_table[395] = 10'h2_08; action_table[396] = 10'h0_00; action_table[397] = 10'h0_00; action_table[398] = 10'h0_00; action_table[399] = 10'h0_00;
action_table[400] = 10'h0_00; action_table[401] = 10'h0_00; action_table[402] = 10'h0_00; action_table[403] = 10'h0_00; action_table[404] = 10'h0_00; action_table[405] = 10'h0_00; action_table[406] = 10'h0_00; action_table[407] = 10'h0_00; action_table[408] = 10'h0_00; action_table[409] = 10'h2_09; action_table[410] = 10'h2_09; action_table[411] = 10'h2_09; action_table[412] = 10'h0_00; action_table[413] = 10'h0_00; action_table[414] = 10'h0_00; action_table[415] = 10'h0_00;
action_table[416] = 10'h2_03; action_table[417] = 10'h2_03; action_table[418] = 10'h2_03; action_table[419] = 10'h0_00; action_table[420] = 10'h2_03; action_table[421] = 10'h2_03; action_table[422] = 10'h2_03; action_table[423] = 10'h2_03; action_table[424] = 10'h0_00; action_table[425] = 10'h0_00; action_table[426] = 10'h0_00; action_table[427] = 10'h0_00; action_table[428] = 10'h2_03; action_table[429] = 10'h0_00; action_table[430] = 10'h0_00; action_table[431] = 10'h0_00;
action_table[432] = 10'h0_00; action_table[433] = 10'h0_00; action_table[434] = 10'h0_00; action_table[435] = 10'h0_00; action_table[436] = 10'h0_00; action_table[437] = 10'h0_00; action_table[438] = 10'h0_00; action_table[439] = 10'h0_00; action_table[440] = 10'h0_00; action_table[441] = 10'h1_0d; action_table[442] = 10'h1_0e; action_table[443] = 10'h1_23; action_table[444] = 10'h0_00; action_table[445] = 10'h0_00; action_table[446] = 10'h0_00; action_table[447] = 10'h0_00;
action_table[448] = 10'h0_00; action_table[449] = 10'h0_00; action_table[450] = 10'h0_00; action_table[451] = 10'h0_00; action_table[452] = 10'h0_00; action_table[453] = 10'h0_00; action_table[454] = 10'h0_00; action_table[455] = 10'h0_00; action_table[456] = 10'h0_00; action_table[457] = 10'h1_0d; action_table[458] = 10'h1_0e; action_table[459] = 10'h1_24; action_table[460] = 10'h0_00; action_table[461] = 10'h0_00; action_table[462] = 10'h0_00; action_table[463] = 10'h0_00;
action_table[464] = 10'h0_00; action_table[465] = 10'h0_00; action_table[466] = 10'h0_00; action_table[467] = 10'h0_00; action_table[468] = 10'h0_00; action_table[469] = 10'h0_00; action_table[470] = 10'h0_00; action_table[471] = 10'h0_00; action_table[472] = 10'h0_00; action_table[473] = 10'h1_0d; action_table[474] = 10'h1_0e; action_table[475] = 10'h1_25; action_table[476] = 10'h0_00; action_table[477] = 10'h0_00; action_table[478] = 10'h0_00; action_table[479] = 10'h0_00;
action_table[480] = 10'h0_00; action_table[481] = 10'h0_00; action_table[482] = 10'h0_00; action_table[483] = 10'h0_00; action_table[484] = 10'h0_00; action_table[485] = 10'h0_00; action_table[486] = 10'h0_00; action_table[487] = 10'h0_00; action_table[488] = 10'h1_26; action_table[489] = 10'h1_20; action_table[490] = 10'h1_21; action_table[491] = 10'h0_00; action_table[492] = 10'h0_00; action_table[493] = 10'h0_00; action_table[494] = 10'h0_00; action_table[495] = 10'h0_00;
action_table[496] = 10'h0_00; action_table[497] = 10'h0_00; action_table[498] = 10'h0_00; action_table[499] = 10'h0_00; action_table[500] = 10'h0_00; action_table[501] = 10'h0_00; action_table[502] = 10'h0_00; action_table[503] = 10'h0_00; action_table[504] = 10'h0_00; action_table[505] = 10'h2_0c; action_table[506] = 10'h2_0c; action_table[507] = 10'h2_0c; action_table[508] = 10'h0_00; action_table[509] = 10'h0_00; action_table[510] = 10'h0_00; action_table[511] = 10'h0_00;
action_table[512] = 10'h1_16; action_table[513] = 10'h0_00; action_table[514] = 10'h0_00; action_table[515] = 10'h0_00; action_table[516] = 10'h0_00; action_table[517] = 10'h0_00; action_table[518] = 10'h0_00; action_table[519] = 10'h1_17; action_table[520] = 10'h0_00; action_table[521] = 10'h0_00; action_table[522] = 10'h0_00; action_table[523] = 10'h0_00; action_table[524] = 10'h0_00; action_table[525] = 10'h0_00; action_table[526] = 10'h0_00; action_table[527] = 10'h0_00;
action_table[528] = 10'h1_16; action_table[529] = 10'h0_00; action_table[530] = 10'h0_00; action_table[531] = 10'h0_00; action_table[532] = 10'h0_00; action_table[533] = 10'h0_00; action_table[534] = 10'h0_00; action_table[535] = 10'h1_17; action_table[536] = 10'h0_00; action_table[537] = 10'h0_00; action_table[538] = 10'h0_00; action_table[539] = 10'h0_00; action_table[540] = 10'h0_00; action_table[541] = 10'h0_00; action_table[542] = 10'h0_00; action_table[543] = 10'h0_00;
action_table[544] = 10'h0_00; action_table[545] = 10'h0_00; action_table[546] = 10'h0_00; action_table[547] = 10'h0_00; action_table[548] = 10'h0_00; action_table[549] = 10'h0_00; action_table[550] = 10'h0_00; action_table[551] = 10'h0_00; action_table[552] = 10'h1_29; action_table[553] = 10'h1_2a; action_table[554] = 10'h1_2b; action_table[555] = 10'h0_00; action_table[556] = 10'h0_00; action_table[557] = 10'h0_00; action_table[558] = 10'h0_00; action_table[559] = 10'h0_00;
action_table[560] = 10'h2_04; action_table[561] = 10'h2_04; action_table[562] = 10'h2_04; action_table[563] = 10'h0_00; action_table[564] = 10'h2_04; action_table[565] = 10'h2_04; action_table[566] = 10'h2_04; action_table[567] = 10'h2_04; action_table[568] = 10'h0_00; action_table[569] = 10'h0_00; action_table[570] = 10'h0_00; action_table[571] = 10'h0_00; action_table[572] = 10'h2_04; action_table[573] = 10'h0_00; action_table[574] = 10'h0_00; action_table[575] = 10'h0_00;
action_table[576] = 10'h2_05; action_table[577] = 10'h2_05; action_table[578] = 10'h2_05; action_table[579] = 10'h0_00; action_table[580] = 10'h2_05; action_table[581] = 10'h2_05; action_table[582] = 10'h2_05; action_table[583] = 10'h2_05; action_table[584] = 10'h0_00; action_table[585] = 10'h0_00; action_table[586] = 10'h0_00; action_table[587] = 10'h0_00; action_table[588] = 10'h2_05; action_table[589] = 10'h0_00; action_table[590] = 10'h0_00; action_table[591] = 10'h0_00;
action_table[592] = 10'h2_06; action_table[593] = 10'h2_06; action_table[594] = 10'h2_06; action_table[595] = 10'h0_00; action_table[596] = 10'h2_06; action_table[597] = 10'h2_06; action_table[598] = 10'h2_06; action_table[599] = 10'h2_06; action_table[600] = 10'h0_00; action_table[601] = 10'h0_00; action_table[602] = 10'h0_00; action_table[603] = 10'h0_00; action_table[604] = 10'h2_06; action_table[605] = 10'h0_00; action_table[606] = 10'h0_00; action_table[607] = 10'h0_00;
action_table[608] = 10'h1_09; action_table[609] = 10'h1_03; action_table[610] = 10'h1_04; action_table[611] = 10'h0_00; action_table[612] = 10'h1_05; action_table[613] = 10'h1_06; action_table[614] = 10'h1_07; action_table[615] = 10'h1_0a; action_table[616] = 10'h0_00; action_table[617] = 10'h0_00; action_table[618] = 10'h0_00; action_table[619] = 10'h0_00; action_table[620] = 10'h0_00; action_table[621] = 10'h0_00; action_table[622] = 10'h0_00; action_table[623] = 10'h0_00;
action_table[624] = 10'h0_00; action_table[625] = 10'h0_00; action_table[626] = 10'h0_00; action_table[627] = 10'h0_00; action_table[628] = 10'h0_00; action_table[629] = 10'h0_00; action_table[630] = 10'h0_00; action_table[631] = 10'h0_00; action_table[632] = 10'h2_08; action_table[633] = 10'h2_08; action_table[634] = 10'h2_08; action_table[635] = 10'h0_00; action_table[636] = 10'h0_00; action_table[637] = 10'h0_00; action_table[638] = 10'h0_00; action_table[639] = 10'h0_00;
action_table[640] = 10'h0_00; action_table[641] = 10'h0_00; action_table[642] = 10'h0_00; action_table[643] = 10'h0_00; action_table[644] = 10'h0_00; action_table[645] = 10'h0_00; action_table[646] = 10'h0_00; action_table[647] = 10'h0_00; action_table[648] = 10'h2_09; action_table[649] = 10'h2_09; action_table[650] = 10'h2_09; action_table[651] = 10'h0_00; action_table[652] = 10'h0_00; action_table[653] = 10'h0_00; action_table[654] = 10'h0_00; action_table[655] = 10'h0_00;
action_table[656] = 10'h0_00; action_table[657] = 10'h0_00; action_table[658] = 10'h0_00; action_table[659] = 10'h0_00; action_table[660] = 10'h0_00; action_table[661] = 10'h0_00; action_table[662] = 10'h0_00; action_table[663] = 10'h0_00; action_table[664] = 10'h2_0c; action_table[665] = 10'h2_0c; action_table[666] = 10'h2_0c; action_table[667] = 10'h0_00; action_table[668] = 10'h0_00; action_table[669] = 10'h0_00; action_table[670] = 10'h0_00; action_table[671] = 10'h0_00;
action_table[672] = 10'h2_07; action_table[673] = 10'h2_07; action_table[674] = 10'h2_07; action_table[675] = 10'h0_00; action_table[676] = 10'h2_07; action_table[677] = 10'h2_07; action_table[678] = 10'h2_07; action_table[679] = 10'h2_07; action_table[680] = 10'h0_00; action_table[681] = 10'h0_00; action_table[682] = 10'h0_00; action_table[683] = 10'h0_00; action_table[684] = 10'h2_07; action_table[685] = 10'h0_00; action_table[686] = 10'h0_00; action_table[687] = 10'h0_00;

reduce_table[0] = 8'h02;
reduce_table[1] = 8'h00;
reduce_table[2] = 8'h02;
reduce_table[3] = 8'h03;
reduce_table[4] = 8'h04;
reduce_table[5] = 8'h04;
reduce_table[6] = 8'h04;
reduce_table[7] = 8'h05;
reduce_table[8] = 8'h03;
reduce_table[9] = 8'h03;
reduce_table[10] = 8'h01;
reduce_table[11] = 8'h01;
reduce_table[12] = 8'h03;

goto_table[0] = 8'h00; goto_table[1] = 8'h00; goto_table[2] = 8'h01; goto_table[3] = 8'h01; goto_table[4] = 8'h01; goto_table[5] = 8'h01; goto_table[6] = 8'h01; goto_table[7] = 8'h01; goto_table[8] = 8'h02; goto_table[9] = 8'h02; goto_table[10] = 8'h02; goto_table[11] = 8'h08; goto_table[12] = 8'h08; goto_table[13] = 8'h00; goto_table[14] = 8'h00; goto_table[15] = 8'h00;
goto_table[16] = 8'h0b; goto_table[17] = 8'h0b; goto_table[18] = 8'h01; goto_table[19] = 8'h01; goto_table[20] = 8'h01; goto_table[21] = 8'h01; goto_table[22] = 8'h01; goto_table[23] = 8'h01; goto_table[24] = 8'h02; goto_table[25] = 8'h02; goto_table[26] = 8'h02; goto_table[27] = 8'h08; goto_table[28] = 8'h08; goto_table[29] = 8'h00; goto_table[30] = 8'h00; goto_table[31] = 8'h00;
goto_table[32] = 8'h00; goto_table[33] = 8'h00; goto_table[34] = 8'h00; goto_table[35] = 8'h00; goto_table[36] = 8'h00; goto_table[37] = 8'h00; goto_table[38] = 8'h00; goto_table[39] = 8'h00; goto_table[40] = 8'h00; goto_table[41] = 8'h00; goto_table[42] = 8'h00; goto_table[43] = 8'h00; goto_table[44] = 8'h00; goto_table[45] = 8'h00; goto_table[46] = 8'h00; goto_table[47] = 8'h00;
goto_table[48] = 8'h00; goto_table[49] = 8'h00; goto_table[50] = 8'h00; goto_table[51] = 8'h00; goto_table[52] = 8'h00; goto_table[53] = 8'h00; goto_table[54] = 8'h00; goto_table[55] = 8'h00; goto_table[56] = 8'h0f; goto_table[57] = 8'h0f; goto_table[58] = 8'h0f; goto_table[59] = 8'h08; goto_table[60] = 8'h08; goto_table[61] = 8'h00; goto_table[62] = 8'h00; goto_table[63] = 8'h00;
goto_table[64] = 8'h00; goto_table[65] = 8'h00; goto_table[66] = 8'h00; goto_table[67] = 8'h00; goto_table[68] = 8'h00; goto_table[69] = 8'h00; goto_table[70] = 8'h00; goto_table[71] = 8'h00; goto_table[72] = 8'h00; goto_table[73] = 8'h00; goto_table[74] = 8'h00; goto_table[75] = 8'h00; goto_table[76] = 8'h00; goto_table[77] = 8'h00; goto_table[78] = 8'h00; goto_table[79] = 8'h00;
goto_table[80] = 8'h00; goto_table[81] = 8'h00; goto_table[82] = 8'h00; goto_table[83] = 8'h00; goto_table[84] = 8'h00; goto_table[85] = 8'h00; goto_table[86] = 8'h00; goto_table[87] = 8'h00; goto_table[88] = 8'h00; goto_table[89] = 8'h00; goto_table[90] = 8'h00; goto_table[91] = 8'h00; goto_table[92] = 8'h00; goto_table[93] = 8'h00; goto_table[94] = 8'h00; goto_table[95] = 8'h00;
goto_table[96] = 8'h00; goto_table[97] = 8'h00; goto_table[98] = 8'h00; goto_table[99] = 8'h00; goto_table[100] = 8'h00; goto_table[101] = 8'h00; goto_table[102] = 8'h00; goto_table[103] = 8'h00; goto_table[104] = 8'h00; goto_table[105] = 8'h00; goto_table[106] = 8'h00; goto_table[107] = 8'h00; goto_table[108] = 8'h00; goto_table[109] = 8'h00; goto_table[110] = 8'h00; goto_table[111] = 8'h00;
goto_table[112] = 8'h00; goto_table[113] = 8'h00; goto_table[114] = 8'h00; goto_table[115] = 8'h00; goto_table[116] = 8'h00; goto_table[117] = 8'h00; goto_table[118] = 8'h00; goto_table[119] = 8'h00; goto_table[120] = 8'h00; goto_table[121] = 8'h00; goto_table[122] = 8'h00; goto_table[123] = 8'h00; goto_table[124] = 8'h00; goto_table[125] = 8'h00; goto_table[126] = 8'h00; goto_table[127] = 8'h00;
goto_table[128] = 8'h00; goto_table[129] = 8'h00; goto_table[130] = 8'h00; goto_table[131] = 8'h00; goto_table[132] = 8'h00; goto_table[133] = 8'h00; goto_table[134] = 8'h00; goto_table[135] = 8'h00; goto_table[136] = 8'h00; goto_table[137] = 8'h00; goto_table[138] = 8'h00; goto_table[139] = 8'h00; goto_table[140] = 8'h00; goto_table[141] = 8'h00; goto_table[142] = 8'h00; goto_table[143] = 8'h00;
goto_table[144] = 8'h00; goto_table[145] = 8'h00; goto_table[146] = 8'h00; goto_table[147] = 8'h00; goto_table[148] = 8'h00; goto_table[149] = 8'h00; goto_table[150] = 8'h00; goto_table[151] = 8'h00; goto_table[152] = 8'h00; goto_table[153] = 8'h00; goto_table[154] = 8'h00; goto_table[155] = 8'h00; goto_table[156] = 8'h00; goto_table[157] = 8'h00; goto_table[158] = 8'h00; goto_table[159] = 8'h00;
goto_table[160] = 8'h00; goto_table[161] = 8'h00; goto_table[162] = 8'h00; goto_table[163] = 8'h00; goto_table[164] = 8'h00; goto_table[165] = 8'h00; goto_table[166] = 8'h00; goto_table[167] = 8'h00; goto_table[168] = 8'h14; goto_table[169] = 8'h14; goto_table[170] = 8'h14; goto_table[171] = 8'h15; goto_table[172] = 8'h15; goto_table[173] = 8'h00; goto_table[174] = 8'h00; goto_table[175] = 8'h00;
goto_table[176] = 8'h00; goto_table[177] = 8'h00; goto_table[178] = 8'h00; goto_table[179] = 8'h00; goto_table[180] = 8'h00; goto_table[181] = 8'h00; goto_table[182] = 8'h00; goto_table[183] = 8'h00; goto_table[184] = 8'h00; goto_table[185] = 8'h00; goto_table[186] = 8'h00; goto_table[187] = 8'h00; goto_table[188] = 8'h00; goto_table[189] = 8'h00; goto_table[190] = 8'h00; goto_table[191] = 8'h00;
goto_table[192] = 8'h00; goto_table[193] = 8'h00; goto_table[194] = 8'h00; goto_table[195] = 8'h00; goto_table[196] = 8'h00; goto_table[197] = 8'h00; goto_table[198] = 8'h00; goto_table[199] = 8'h00; goto_table[200] = 8'h00; goto_table[201] = 8'h00; goto_table[202] = 8'h00; goto_table[203] = 8'h00; goto_table[204] = 8'h00; goto_table[205] = 8'h00; goto_table[206] = 8'h00; goto_table[207] = 8'h00;
goto_table[208] = 8'h00; goto_table[209] = 8'h00; goto_table[210] = 8'h00; goto_table[211] = 8'h00; goto_table[212] = 8'h00; goto_table[213] = 8'h00; goto_table[214] = 8'h00; goto_table[215] = 8'h00; goto_table[216] = 8'h00; goto_table[217] = 8'h00; goto_table[218] = 8'h00; goto_table[219] = 8'h18; goto_table[220] = 8'h18; goto_table[221] = 8'h00; goto_table[222] = 8'h00; goto_table[223] = 8'h00;
goto_table[224] = 8'h00; goto_table[225] = 8'h00; goto_table[226] = 8'h00; goto_table[227] = 8'h00; goto_table[228] = 8'h00; goto_table[229] = 8'h00; goto_table[230] = 8'h00; goto_table[231] = 8'h00; goto_table[232] = 8'h00; goto_table[233] = 8'h00; goto_table[234] = 8'h00; goto_table[235] = 8'h19; goto_table[236] = 8'h19; goto_table[237] = 8'h00; goto_table[238] = 8'h00; goto_table[239] = 8'h00;
goto_table[240] = 8'h00; goto_table[241] = 8'h00; goto_table[242] = 8'h00; goto_table[243] = 8'h00; goto_table[244] = 8'h00; goto_table[245] = 8'h00; goto_table[246] = 8'h00; goto_table[247] = 8'h00; goto_table[248] = 8'h00; goto_table[249] = 8'h00; goto_table[250] = 8'h00; goto_table[251] = 8'h00; goto_table[252] = 8'h00; goto_table[253] = 8'h00; goto_table[254] = 8'h00; goto_table[255] = 8'h00;
goto_table[256] = 8'h00; goto_table[257] = 8'h00; goto_table[258] = 8'h00; goto_table[259] = 8'h00; goto_table[260] = 8'h00; goto_table[261] = 8'h00; goto_table[262] = 8'h00; goto_table[263] = 8'h00; goto_table[264] = 8'h1b; goto_table[265] = 8'h1b; goto_table[266] = 8'h1b; goto_table[267] = 8'h08; goto_table[268] = 8'h08; goto_table[269] = 8'h00; goto_table[270] = 8'h00; goto_table[271] = 8'h00;
goto_table[272] = 8'h00; goto_table[273] = 8'h00; goto_table[274] = 8'h00; goto_table[275] = 8'h00; goto_table[276] = 8'h00; goto_table[277] = 8'h00; goto_table[278] = 8'h00; goto_table[279] = 8'h00; goto_table[280] = 8'h1c; goto_table[281] = 8'h1c; goto_table[282] = 8'h1c; goto_table[283] = 8'h08; goto_table[284] = 8'h08; goto_table[285] = 8'h00; goto_table[286] = 8'h00; goto_table[287] = 8'h00;
goto_table[288] = 8'h00; goto_table[289] = 8'h00; goto_table[290] = 8'h00; goto_table[291] = 8'h00; goto_table[292] = 8'h00; goto_table[293] = 8'h00; goto_table[294] = 8'h00; goto_table[295] = 8'h00; goto_table[296] = 8'h1d; goto_table[297] = 8'h1d; goto_table[298] = 8'h1d; goto_table[299] = 8'h08; goto_table[300] = 8'h08; goto_table[301] = 8'h00; goto_table[302] = 8'h00; goto_table[303] = 8'h00;
goto_table[304] = 8'h00; goto_table[305] = 8'h00; goto_table[306] = 8'h00; goto_table[307] = 8'h00; goto_table[308] = 8'h00; goto_table[309] = 8'h00; goto_table[310] = 8'h00; goto_table[311] = 8'h00; goto_table[312] = 8'h1e; goto_table[313] = 8'h1e; goto_table[314] = 8'h1e; goto_table[315] = 8'h15; goto_table[316] = 8'h15; goto_table[317] = 8'h00; goto_table[318] = 8'h00; goto_table[319] = 8'h00;
goto_table[320] = 8'h00; goto_table[321] = 8'h00; goto_table[322] = 8'h00; goto_table[323] = 8'h00; goto_table[324] = 8'h00; goto_table[325] = 8'h00; goto_table[326] = 8'h00; goto_table[327] = 8'h00; goto_table[328] = 8'h00; goto_table[329] = 8'h00; goto_table[330] = 8'h00; goto_table[331] = 8'h00; goto_table[332] = 8'h00; goto_table[333] = 8'h00; goto_table[334] = 8'h00; goto_table[335] = 8'h00;
goto_table[336] = 8'h00; goto_table[337] = 8'h00; goto_table[338] = 8'h00; goto_table[339] = 8'h00; goto_table[340] = 8'h00; goto_table[341] = 8'h00; goto_table[342] = 8'h00; goto_table[343] = 8'h00; goto_table[344] = 8'h00; goto_table[345] = 8'h00; goto_table[346] = 8'h00; goto_table[347] = 8'h00; goto_table[348] = 8'h00; goto_table[349] = 8'h00; goto_table[350] = 8'h00; goto_table[351] = 8'h00;
goto_table[352] = 8'h00; goto_table[353] = 8'h00; goto_table[354] = 8'h00; goto_table[355] = 8'h00; goto_table[356] = 8'h00; goto_table[357] = 8'h00; goto_table[358] = 8'h00; goto_table[359] = 8'h00; goto_table[360] = 8'h00; goto_table[361] = 8'h00; goto_table[362] = 8'h00; goto_table[363] = 8'h00; goto_table[364] = 8'h00; goto_table[365] = 8'h00; goto_table[366] = 8'h00; goto_table[367] = 8'h00;
goto_table[368] = 8'h00; goto_table[369] = 8'h00; goto_table[370] = 8'h00; goto_table[371] = 8'h00; goto_table[372] = 8'h00; goto_table[373] = 8'h00; goto_table[374] = 8'h00; goto_table[375] = 8'h00; goto_table[376] = 8'h22; goto_table[377] = 8'h22; goto_table[378] = 8'h22; goto_table[379] = 8'h15; goto_table[380] = 8'h15; goto_table[381] = 8'h00; goto_table[382] = 8'h00; goto_table[383] = 8'h00;
goto_table[384] = 8'h00; goto_table[385] = 8'h00; goto_table[386] = 8'h00; goto_table[387] = 8'h00; goto_table[388] = 8'h00; goto_table[389] = 8'h00; goto_table[390] = 8'h00; goto_table[391] = 8'h00; goto_table[392] = 8'h00; goto_table[393] = 8'h00; goto_table[394] = 8'h00; goto_table[395] = 8'h00; goto_table[396] = 8'h00; goto_table[397] = 8'h00; goto_table[398] = 8'h00; goto_table[399] = 8'h00;
goto_table[400] = 8'h00; goto_table[401] = 8'h00; goto_table[402] = 8'h00; goto_table[403] = 8'h00; goto_table[404] = 8'h00; goto_table[405] = 8'h00; goto_table[406] = 8'h00; goto_table[407] = 8'h00; goto_table[408] = 8'h00; goto_table[409] = 8'h00; goto_table[410] = 8'h00; goto_table[411] = 8'h00; goto_table[412] = 8'h00; goto_table[413] = 8'h00; goto_table[414] = 8'h00; goto_table[415] = 8'h00;
goto_table[416] = 8'h00; goto_table[417] = 8'h00; goto_table[418] = 8'h00; goto_table[419] = 8'h00; goto_table[420] = 8'h00; goto_table[421] = 8'h00; goto_table[422] = 8'h00; goto_table[423] = 8'h00; goto_table[424] = 8'h00; goto_table[425] = 8'h00; goto_table[426] = 8'h00; goto_table[427] = 8'h00; goto_table[428] = 8'h00; goto_table[429] = 8'h00; goto_table[430] = 8'h00; goto_table[431] = 8'h00;
goto_table[432] = 8'h00; goto_table[433] = 8'h00; goto_table[434] = 8'h00; goto_table[435] = 8'h00; goto_table[436] = 8'h00; goto_table[437] = 8'h00; goto_table[438] = 8'h00; goto_table[439] = 8'h00; goto_table[440] = 8'h00; goto_table[441] = 8'h00; goto_table[442] = 8'h00; goto_table[443] = 8'h00; goto_table[444] = 8'h00; goto_table[445] = 8'h00; goto_table[446] = 8'h00; goto_table[447] = 8'h00;
goto_table[448] = 8'h00; goto_table[449] = 8'h00; goto_table[450] = 8'h00; goto_table[451] = 8'h00; goto_table[452] = 8'h00; goto_table[453] = 8'h00; goto_table[454] = 8'h00; goto_table[455] = 8'h00; goto_table[456] = 8'h00; goto_table[457] = 8'h00; goto_table[458] = 8'h00; goto_table[459] = 8'h00; goto_table[460] = 8'h00; goto_table[461] = 8'h00; goto_table[462] = 8'h00; goto_table[463] = 8'h00;
goto_table[464] = 8'h00; goto_table[465] = 8'h00; goto_table[466] = 8'h00; goto_table[467] = 8'h00; goto_table[468] = 8'h00; goto_table[469] = 8'h00; goto_table[470] = 8'h00; goto_table[471] = 8'h00; goto_table[472] = 8'h00; goto_table[473] = 8'h00; goto_table[474] = 8'h00; goto_table[475] = 8'h00; goto_table[476] = 8'h00; goto_table[477] = 8'h00; goto_table[478] = 8'h00; goto_table[479] = 8'h00;
goto_table[480] = 8'h00; goto_table[481] = 8'h00; goto_table[482] = 8'h00; goto_table[483] = 8'h00; goto_table[484] = 8'h00; goto_table[485] = 8'h00; goto_table[486] = 8'h00; goto_table[487] = 8'h00; goto_table[488] = 8'h00; goto_table[489] = 8'h00; goto_table[490] = 8'h00; goto_table[491] = 8'h00; goto_table[492] = 8'h00; goto_table[493] = 8'h00; goto_table[494] = 8'h00; goto_table[495] = 8'h00;
goto_table[496] = 8'h00; goto_table[497] = 8'h00; goto_table[498] = 8'h00; goto_table[499] = 8'h00; goto_table[500] = 8'h00; goto_table[501] = 8'h00; goto_table[502] = 8'h00; goto_table[503] = 8'h00; goto_table[504] = 8'h00; goto_table[505] = 8'h00; goto_table[506] = 8'h00; goto_table[507] = 8'h00; goto_table[508] = 8'h00; goto_table[509] = 8'h00; goto_table[510] = 8'h00; goto_table[511] = 8'h00;
goto_table[512] = 8'h00; goto_table[513] = 8'h00; goto_table[514] = 8'h00; goto_table[515] = 8'h00; goto_table[516] = 8'h00; goto_table[517] = 8'h00; goto_table[518] = 8'h00; goto_table[519] = 8'h00; goto_table[520] = 8'h00; goto_table[521] = 8'h00; goto_table[522] = 8'h00; goto_table[523] = 8'h27; goto_table[524] = 8'h27; goto_table[525] = 8'h00; goto_table[526] = 8'h00; goto_table[527] = 8'h00;
goto_table[528] = 8'h00; goto_table[529] = 8'h00; goto_table[530] = 8'h00; goto_table[531] = 8'h00; goto_table[532] = 8'h00; goto_table[533] = 8'h00; goto_table[534] = 8'h00; goto_table[535] = 8'h00; goto_table[536] = 8'h00; goto_table[537] = 8'h00; goto_table[538] = 8'h00; goto_table[539] = 8'h28; goto_table[540] = 8'h28; goto_table[541] = 8'h00; goto_table[542] = 8'h00; goto_table[543] = 8'h00;
goto_table[544] = 8'h00; goto_table[545] = 8'h00; goto_table[546] = 8'h00; goto_table[547] = 8'h00; goto_table[548] = 8'h00; goto_table[549] = 8'h00; goto_table[550] = 8'h00; goto_table[551] = 8'h00; goto_table[552] = 8'h00; goto_table[553] = 8'h00; goto_table[554] = 8'h00; goto_table[555] = 8'h00; goto_table[556] = 8'h00; goto_table[557] = 8'h00; goto_table[558] = 8'h00; goto_table[559] = 8'h00;
goto_table[560] = 8'h00; goto_table[561] = 8'h00; goto_table[562] = 8'h00; goto_table[563] = 8'h00; goto_table[564] = 8'h00; goto_table[565] = 8'h00; goto_table[566] = 8'h00; goto_table[567] = 8'h00; goto_table[568] = 8'h00; goto_table[569] = 8'h00; goto_table[570] = 8'h00; goto_table[571] = 8'h00; goto_table[572] = 8'h00; goto_table[573] = 8'h00; goto_table[574] = 8'h00; goto_table[575] = 8'h00;
goto_table[576] = 8'h00; goto_table[577] = 8'h00; goto_table[578] = 8'h00; goto_table[579] = 8'h00; goto_table[580] = 8'h00; goto_table[581] = 8'h00; goto_table[582] = 8'h00; goto_table[583] = 8'h00; goto_table[584] = 8'h00; goto_table[585] = 8'h00; goto_table[586] = 8'h00; goto_table[587] = 8'h00; goto_table[588] = 8'h00; goto_table[589] = 8'h00; goto_table[590] = 8'h00; goto_table[591] = 8'h00;
goto_table[592] = 8'h00; goto_table[593] = 8'h00; goto_table[594] = 8'h00; goto_table[595] = 8'h00; goto_table[596] = 8'h00; goto_table[597] = 8'h00; goto_table[598] = 8'h00; goto_table[599] = 8'h00; goto_table[600] = 8'h00; goto_table[601] = 8'h00; goto_table[602] = 8'h00; goto_table[603] = 8'h00; goto_table[604] = 8'h00; goto_table[605] = 8'h00; goto_table[606] = 8'h00; goto_table[607] = 8'h00;
goto_table[608] = 8'h00; goto_table[609] = 8'h00; goto_table[610] = 8'h2a; goto_table[611] = 8'h2a; goto_table[612] = 8'h2a; goto_table[613] = 8'h2a; goto_table[614] = 8'h2a; goto_table[615] = 8'h2a; goto_table[616] = 8'h02; goto_table[617] = 8'h02; goto_table[618] = 8'h02; goto_table[619] = 8'h08; goto_table[620] = 8'h08; goto_table[621] = 8'h00; goto_table[622] = 8'h00; goto_table[623] = 8'h00;
goto_table[624] = 8'h00; goto_table[625] = 8'h00; goto_table[626] = 8'h00; goto_table[627] = 8'h00; goto_table[628] = 8'h00; goto_table[629] = 8'h00; goto_table[630] = 8'h00; goto_table[631] = 8'h00; goto_table[632] = 8'h00; goto_table[633] = 8'h00; goto_table[634] = 8'h00; goto_table[635] = 8'h00; goto_table[636] = 8'h00; goto_table[637] = 8'h00; goto_table[638] = 8'h00; goto_table[639] = 8'h00;
goto_table[640] = 8'h00; goto_table[641] = 8'h00; goto_table[642] = 8'h00; goto_table[643] = 8'h00; goto_table[644] = 8'h00; goto_table[645] = 8'h00; goto_table[646] = 8'h00; goto_table[647] = 8'h00; goto_table[648] = 8'h00; goto_table[649] = 8'h00; goto_table[650] = 8'h00; goto_table[651] = 8'h00; goto_table[652] = 8'h00; goto_table[653] = 8'h00; goto_table[654] = 8'h00; goto_table[655] = 8'h00;
goto_table[656] = 8'h00; goto_table[657] = 8'h00; goto_table[658] = 8'h00; goto_table[659] = 8'h00; goto_table[660] = 8'h00; goto_table[661] = 8'h00; goto_table[662] = 8'h00; goto_table[663] = 8'h00; goto_table[664] = 8'h00; goto_table[665] = 8'h00; goto_table[666] = 8'h00; goto_table[667] = 8'h00; goto_table[668] = 8'h00; goto_table[669] = 8'h00; goto_table[670] = 8'h00; goto_table[671] = 8'h00;
goto_table[672] = 8'h00; goto_table[673] = 8'h00; goto_table[674] = 8'h00; goto_table[675] = 8'h00; goto_table[676] = 8'h00; goto_table[677] = 8'h00; goto_table[678] = 8'h00; goto_table[679] = 8'h00; goto_table[680] = 8'h00; goto_table[681] = 8'h00; goto_table[682] = 8'h00; goto_table[683] = 8'h00; goto_table[684] = 8'h00; goto_table[685] = 8'h00; goto_table[686] = 8'h00; goto_table[687] = 8'h00;
